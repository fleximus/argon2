module argon2

fn test_simple_argon2i() {
	result := hash_i_raw(2, 65536, 1, 'password'.bytes(), 'somesalt'.bytes(), 32) or { panic(err) }
	expected := [u8(0xc1), 0x62, 0x88, 0x32, 0x14, 0x7d, 0x97, 0x20, 0xc5, 0xbd, 0x1c, 0xfd, 0x61, 0x36, 0x70, 0x78, 0x72, 0x9f, 0x6d, 0xfb, 0x6f, 0x8f, 0xea, 0x9f, 0xf9, 0x81, 0x58, 0xe0, 0xd7, 0x81, 0x6e, 0xd0]
	
	
	assert result == expected, 'Argon2i test should match expected hash'
}

